netcdf depth_axis_test {
dimensions:
	depth_p1 = 31 ;
	depth = 30 ;
variables:
	double depth_edges(depth_p1) ;
		depth_edges:long_name = "Depth Layer Edges" ;
		depth_edges:units = "m" ;
	double depth_delta(depth) ;
		depth_delta:long_name = "Depth Layer Thickness" ;
		depth_delta:units = "m" ;
data:

 depth_edges = 0, 10, 20, 30, 40, 50, 60, 70, 80, 92, 106, 122, 140, 160, 
    182, 206, 232, 260, 290, 320, 350, 380, 410, 440, 470, 500, 530, 560, 
    590, 620, 650 ;

 depth_delta = 10, 10, 10, 10, 10, 10, 10, 10, 12, 14, 16, 18, 20, 22, 24, 
    26, 28, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30 ;
}
